module tb(
input wreq,rreq,
input clk,
input  [7:0] wdata,
input rst,
output  [7:0] rdata;
output f,e

);

endmodule